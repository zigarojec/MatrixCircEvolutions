* wrapping circuit for arithmetic circuit evolution
* Ziga Rojec, EDA, FE, UL, 2021

*.include 'models_for_start.inc'
*.include 'rectifier.cir'

xcirc vin inb vout 0 HOT_CIRCUIT

*****Power supply*****
*vdd (vdd 0) dc = 12

******Input resistors*****
*r0    (vin vout) r=10k

vin (vin inb) dc = 10

*****Loads*****
*.param rl=1000k
*rl (vout 0) r=1meg
*rl (vout 0) r=1k
rl (vout voutm) r=1k
vl (voutm 0) dc=0


*.end
