
.subckt 