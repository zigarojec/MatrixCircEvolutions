* wrapping circuit for arithmetic circuit evolution
* Ziga Rojec, EDA, FE, UL, 2021


*.include 'models_for_start.inc'
*.include 'scoreCirc_squareroot_resilenceMode_g_0_i_0_subckt.cir'

xcirc vout 0 HOT_CIRCUIT

*****Power supply*****
*vdd (vdd 0) dc = 12

******Input resistors*****
r0    (vin vout) r=10k

vin (vin 0) dc = 10

*****Loads*****
*.param rl=1000k
rl (vout 0) r=1meg


*.end
